* C:\LTSpiceTransmissionLines\LTSpice\sim\main\tranmission_line_14_dropoffs.asc
O2 N014 N028 Out OutRef LossyTL
rf N028 0 100k
C1 N014 0 {Cdrp}
O1 N013 N027 N014 N028 LossyTL
rf1 N027 0 100k
C2 N013 0 {Cdrp}
O3 N012 N026 N013 N027 LossyTL
rf2 N026 0 100k
C3 N012 0 {Cdrp}
O4 N011 N025 N012 N026 LossyTL
rf3 N025 0 100k
C4 N011 0 {Cdrp}
O5 N010 N024 N011 N025 LossyTL
rf4 N024 0 100k
C5 N010 0 {Cdrp}
O6 N009 N023 N010 N024 LossyTL
rf5 N023 0 100k
C6 N009 0 {Cdrp}
O7 N008 N022 N009 N023 LossyTL
rf6 N022 0 100k
C7 N008 0 {Cdrp}
O8 N007 N021 N008 N022 LossyTL
rf7 N021 0 100k
C8 N007 0 {Cdrp}
O9 N006 N020 N007 N021 LossyTL
rf8 N020 0 100k
C9 N006 0 {Cdrp}
O10 N005 N019 N006 N020 LossyTL
rf9 N019 0 100k
C10 N005 0 {Cdrp}
O11 N004 N018 N005 N019 LossyTL
rf10 N018 0 100k
C11 N004 0 {Cdrp}
O12 N003 N017 N004 N018 LossyTL
rf11 N017 0 100k
C12 N003 0 {Cdrp}
O13 N002 N016 N003 N017 LossyTL
rf12 N016 0 100k
C13 N002 0 {Cdrp}
O14 N001 N015 N002 N016 LossyTL
rf13 N015 0 100k
C14 N001 0 {Cdrp}
RoutRef OutRef 0 100k
O27 InPulse InRefPulse N001 N015 LossyTL
R16 InPulse InRefPulse {Rterm}
R17 InRefPulse 0 100k
V2 InPulse InRefPulse PULSE(0 1 0 2n 2n 16n) AC 1 Rser=0
R2 Out OutRef {Rterm}
.model LossyTL  LTRA(len=Lenline R=Rline L=Lline C=Cline)
.tran 0 100n
;ac oct 50 10k 1000Meg
;step param Rline 0.02 2 0.2
;step param Lline 0.079n 7.9n 0.79n
;step param Cline 0.22p 22p 2.2p
;step param Cdrp 1p 5p 1p
;step param Lenline 1.0 10.0 1.0
.param  Cdrp = 1p  Rterm =sqrt(Lline/Cline) Lenline=5 Rline=1.02 Lline=1.659n Cline=2.42p
.save V(Out) V(N001) V(N015) V(N014) V(N028) V(N008) V(N022) V(InPulse)
.backanno
.end
