* C:\LTSpiceTransmissionLines\LTSpice\sim\main\tranmission_line_10_dropoffs.asc
O2 N010 N020 Out OutRef LossyTL
rf N020 0 100k
C1 N010 N020 {Cdrp}
O1 N009 N019 N010 N020 LossyTL
rf1 N019 0 100k
C2 N009 N019 {Cdrp}
O3 N008 N018 N009 N019 LossyTL
rf2 N018 0 100k
C3 N008 N018 {Cdrp}
O4 N007 N017 N008 N018 LossyTL
rf3 N017 0 100k
C4 N007 N017 {Cdrp}
O5 N006 N016 N007 N017 LossyTL
rf4 N016 0 100k
C5 N006 N016 {Cdrp}
O6 N005 N015 N006 N016 LossyTL
rf5 N015 0 100k
C6 N005 N015 {Cdrp}
O7 N004 N014 N005 N015 LossyTL
rf6 N014 0 100k
C7 N004 N014 {Cdrp}
O8 N003 N013 N004 N014 LossyTL
rf7 N013 0 100k
C8 N003 N013 {Cdrp}
O9 N002 N012 N003 N013 LossyTL
rf8 N012 0 100k
C9 N002 N012 {Cdrp}
O10 N001 N011 N002 N012 LossyTL
rf9 N011 0 100k
C10 N001 N011 {Cdrp}
RoutRef OutRef 0 100k
O27 InPulse InRefPulse N001 N011 LossyTL
R16 InPulse InRefPulse {Rterm}
R17 InRefPulse 0 100k
R2 Out OutRef {Rterm}
I1 InPulse InRefPulse PULSE(0 -50m 0 100p 100p 1.5n) AC 1
I2 InPulse InRefPulse PULSE(0 0 1.5n 100p 100p 1.3n) AC 1
I3 InPulse InRefPulse PULSE(0 -50m 3n 100p 100p 1.3n) AC 1
I4 InPulse InRefPulse PULSE(0 0 4.5n 100p 100p 1.3n) AC 1
I5 InPulse InRefPulse PULSE(0 -50m 6n 100p 100p 1.3n) AC 1
.tran 0 100n
;ac oct 50 10k 1000Meg
;step param Rline 0.02 2 .8
;step param Lline 0.079n 7.9n 3.16n
;step param Cline 0.22p 22p 8.8p
.param  Cdrp = 1p  Rterm =sqrt(Lline/Cline) Lenline=5 Rline=1.02 Lline=1.659n Cline=2.42p
.save V(Out) V(N001) V(N010) V(N006) V(InPulse)
.model LossyTL  LTRA(len=Lenline R=Rline L=Lline C=Cline)
.backanno
.end
