*5.0pLTSpiceTransmissionLines\LTSpice\sim\main\tranmission_line_10_dropoffs.asc
O2 N010 N020 Out OutRef LossyTL
rf N020 0 100k
C1 N010 0 {Cdrp}
O1 N009 N019 N010 N020 LossyTL
rf1 N019 0 100k
C2 N009 0 {Cdrp}
O3 N008 N018 N009 N019 LossyTL
rf2 N018 0 100k
C3 N008 0 {Cdrp}
O4 N007 N017 N008 N018 LossyTL
rf3 N017 0 100k
C4 N007 0 {Cdrp}
O5 N006 N016 N007 N017 LossyTL
rf4 N016 0 100k
C5 N006 0 {Cdrp}
O6 N005 N015 N006 N016 LossyTL
rf5 N015 0 100k
C6 N005 0 {Cdrp}
O7 N004 N014 N005 N015 LossyTL
rf6 N014 0 100k
C7 N004 0 {Cdrp}
O8 N003 N013 N004 N014 LossyTL
rf7 N013 0 100k
C8 N003 0 {Cdrp}
O9 N002 N012 N003 N013 LossyTL
rf8 N012 0 100k
C9 N002 0 {Cdrp}
O10 N001 N011 N002 N012 LossyTL
rf9 N011 0 100k
C10 N001 0 {Cdrp}
RoutRef OutRef 0 100k
O27 InPulse InRefPulse N001 N011 LossyTL
R16 InPulse InRefPulse {Rterm}
R17 InRefPulse 0 100k
V2 InPulse InRefPulse PULSE(0 1 0 2n 2n 16n) AC 1 Rser=0
R2 Out OutRef {Rterm}
.tran 0 100n
;ac oct 50 10k 1000Meg
;step param Rline 0.02 2 0.2
;step param Lline 0.079n 7.9n 0.79n
;step param Cline 0.22p 22p 2.2p
;step param Cdrp 1p 5p 1p
;step param Lenline 1.0 10.0 1.0
.param  Cdrp=1.0p   Rterm =sqrt(Lline/Cline) Lenline=5.0    Rline=220m  Lline=79.p    Cline=220f
.save V(Out) V(N001) V(N011) V(N010) V(N020) V(N006) V(N016) V(InPulse)
.model LossyTL  LTRA(len=Lenline R=Rline L=Lline C=Cline)
.backanno
.end
